`timescale 1ns/1ns

module WbStage(input clk, input rst);
  
endmodule
