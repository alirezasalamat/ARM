`include "defines.v"

module ExeReg(input clk, input rst);
  
endmodule
