`timescale 1ns/1ns

module IdStage(input clk, input rst);
  
endmodule
