`include "defines.v"

module MemReg(input clk, input rst);
  
endmodule
