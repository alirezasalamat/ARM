`include "defines.v"

module WbStage(input clk, input rst);
  
endmodule
