`include "defines.v"

module IdReg(input clk, input rst);
    
endmodule
