`timescale 1ns/1ns

module test();
  
endmodule
