`timescale 1ns/1ns

module ExeReg(input clk, input rst);
  
endmodule
