`timescale 1ns/1ns

module ExeStage(input clk, input rst);
  
endmodule
