`timescale 1ns/1ns

module IfReg(input clk, input rst);
  
endmodule
