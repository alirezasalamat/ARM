`include "defines.v"

module ExeStage(input clk, input rst);
  
endmodule
