`include "defines.v"

module test();
  
endmodule
