`timescale 1ns/1ns

module IdReg(input clk, input rst);
  
endmodule
