`timescale 1ns/1ns

module MemReg(input clk, input rst);
  
endmodule
