`timescale 1ns/1ns

module MemStage(input clk, input rst);
  
endmodule
