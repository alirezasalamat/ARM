`include "defines.v"

module MemStage(input clk, input rst);
  
endmodule
