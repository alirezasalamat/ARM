`timescale 1ns/1ns

module IfStage(input clk, input rst);
  
endmodule
